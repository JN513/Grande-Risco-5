module mux_tb();

logic [31:0] MUX_A, MUX_B;
logic MUX_Option;
logic [31:0] MUX_S;

MUX MUX(
    .A(MUX_A),
    .B(MUX_B),
    .S(MUX_S),
    .option(MUX_Option)
);

initial begin
    MUX_A = 5;
    MUX_B = 3;
    MUX_Option = 0;

    #1

    $display("Estado ", MUX_S);
    MUX_Option = 1;

    #1
    $display("Estado ", MUX_S);

end

endmodule
