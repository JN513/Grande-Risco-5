module IR_Decompression (
    input wire clk,
    input wire [15:0] compressed_instruction,
    output reg [31:0] decompressed_instruction
);



endmodule