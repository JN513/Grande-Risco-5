`define ENABLE_MDU 1
//`define ENABLE_FPU 1
//`define ENABLE_BMU 1
`define FPGA 1