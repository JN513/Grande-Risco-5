module BMU ( // Bit manipulation unit for riscv B extension
    input wire clk
);
    
endmodule
