module Branch_Prediction (
    input  logic [31:0] PC,
    input  logic [31:0] instruction_data,
    output logic [31:0] address
);
    
endmodule
