module Branch_Prediction (
    input wire [31:0] PC,
    input wire [31:0] instruction_data,
    output wire [31:0] address
);
    
endmodule
